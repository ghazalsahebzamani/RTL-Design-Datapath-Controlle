module merg(input[7:0]p,a,output[15:0]r);
  assign r={p,a};
endmodule

